//`define FASTBOOT
`define SIMULATION