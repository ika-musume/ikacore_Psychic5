/*
    PROM
*/

module PROM #(parameter aw=10, dw=8, pol=1, simhexfile="")
(
    //data loader
    input   wire            i_EMU_PROG_CLK,
    input   wire   [aw-1:0] i_EMU_PROG_ADDR,
    input   wire   [dw-1:0] i_EMU_PROG_DIN,
    input   wire            i_EMU_PROG_CS_n,
    input   wire            i_EMU_PROG_WR_n,
    
    //PCB ports
    input   wire            i_MCLK,
    input   wire   [aw-1:0] i_ADDR,
    output  reg    [dw-1:0] o_DOUT,
    input   wire            i_CS_n,
    input   wire            i_RD_n
);

reg     [dw-1:0]   ROM [0:(2**aw)-1];

generate
    if(pol == 1'b1)
    begin
        always @(posedge i_MCLK) //read
        begin
            if(i_EMU_PROG_CS_n == 1'b1)
            begin
                if(i_CS_n == 1'b0)
                begin
                    if(i_RD_n == 1'b0)
                    begin
                        o_DOUT <= ROM[i_ADDR];
                    end
                end
            end
        end
    end

    else
    begin
        always @(negedge i_MCLK) //read
        begin
            if(i_EMU_PROG_CS_n == 1'b1)
            begin
                if(i_CS_n == 1'b0)
                begin
                    if(i_RD_n == 1'b0)
                    begin
                        o_DOUT <= ROM[i_ADDR];
                    end
                end
            end
        end
    end
endgenerate

always @(posedge i_EMU_PROG_CLK)
begin
    if(i_EMU_PROG_CS_n == 1'b0)
    begin
        if(i_EMU_PROG_WR_n == 1'b0)
        begin
            ROM[i_EMU_PROG_ADDR] <= i_EMU_PROG_DIN;
        end
    end
end

initial
begin
    if( simhexfile != "" ) begin
        $readmemh(simhexfile, ROM);
    end
end

endmodule
